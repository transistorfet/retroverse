module k30logic_tb();

    k30logic DTS(

    );

    

endmodule
